module OneBitCounter
(input clk, input rst, output out)

endmodule 